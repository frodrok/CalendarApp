test.test = Kalender
login = Logga in
register = Registrera dig
username = Användarnamn
password = Lösenord
title = YHC3LKalender